
interface and2_if();

  logic a,b;
  logic c;
endinterface:and2_if


